module fc_rd_ctrl
(
	input clk, rst_n,
