module fc_ctrl
(
	input clk, rst_n,
