module fc_unit
(
	input clk, rst_n,
