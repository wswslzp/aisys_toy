module sys_state_ctrl
(
	// from outside 
	input clk, rst_n,
	
	// uart side
	input 
