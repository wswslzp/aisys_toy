module uart_rd_bridge
(
	input 
